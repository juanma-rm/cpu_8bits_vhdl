----------------------------------------------------------------------------------
----------------------------------------------------------------------------------
-- cpu_octobits.vhd

--! @todo doc
----------------------------------------------------------------------------------
----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
-- Import of libraries and packages
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.utils.all;

----------------------------------------------------------------------------------
-- Entity
----------------------------------------------------------------------------------

entity top is

end top;

----------------------------------------------------------------------------------
-- Architecture
----------------------------------------------------------------------------------

architecture behavioural of top is



begin



end behavioural;
